// nios2_cpu.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module nios2_cpu (
		input  wire        accel_interrupt_export, // accel_interrupt.export
		input  wire [15:0] accel_xdata_export,     //     accel_xdata.export
		input  wire [15:0] accel_ydata_export,     //     accel_ydata.export
		input  wire [15:0] accel_zdata_export,     //     accel_zdata.export
		input  wire        clk_clk,                //             clk.clk
		output wire [7:0]  disp0_export,           //           disp0.export
		output wire [7:0]  disp1_export,           //           disp1.export
		output wire [9:0]  led_export,             //             led.export
		input  wire        reset_reset_n,          //           reset.reset_n
		input  wire [9:0]  switch_export,          //          switch.export
		output wire [8:0]  update_control_export,  //  update_control.export
		output wire [15:0] update_value_export,    //    update_value.export
		output wire [1:0]  x_coeff_bank_export,    //    x_coeff_bank.export
		output wire [1:0]  y_coeff_bank_export,    //    y_coeff_bank.export
		output wire [1:0]  z_coeff_bank_export     //    z_coeff_bank.export
	);

	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [19:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [19:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;          // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;            // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_0_s1_address;             // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;          // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;               // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;           // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;               // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_accel_data_interrupt_s1_chipselect;      // mm_interconnect_0:accel_data_interrupt_s1_chipselect -> accel_data_interrupt:chipselect
	wire  [31:0] mm_interconnect_0_accel_data_interrupt_s1_readdata;        // accel_data_interrupt:readdata -> mm_interconnect_0:accel_data_interrupt_s1_readdata
	wire   [1:0] mm_interconnect_0_accel_data_interrupt_s1_address;         // mm_interconnect_0:accel_data_interrupt_s1_address -> accel_data_interrupt:address
	wire         mm_interconnect_0_accel_data_interrupt_s1_write;           // mm_interconnect_0:accel_data_interrupt_s1_write -> accel_data_interrupt:write_n
	wire  [31:0] mm_interconnect_0_accel_data_interrupt_s1_writedata;       // mm_interconnect_0:accel_data_interrupt_s1_writedata -> accel_data_interrupt:writedata
	wire  [31:0] mm_interconnect_0_accel_xread_s1_readdata;                 // accel_xread:readdata -> mm_interconnect_0:accel_xread_s1_readdata
	wire   [1:0] mm_interconnect_0_accel_xread_s1_address;                  // mm_interconnect_0:accel_xread_s1_address -> accel_xread:address
	wire         mm_interconnect_0_print0_s1_chipselect;                    // mm_interconnect_0:print0_s1_chipselect -> print0:chipselect
	wire  [31:0] mm_interconnect_0_print0_s1_readdata;                      // print0:readdata -> mm_interconnect_0:print0_s1_readdata
	wire   [1:0] mm_interconnect_0_print0_s1_address;                       // mm_interconnect_0:print0_s1_address -> print0:address
	wire         mm_interconnect_0_print0_s1_write;                         // mm_interconnect_0:print0_s1_write -> print0:write_n
	wire  [31:0] mm_interconnect_0_print0_s1_writedata;                     // mm_interconnect_0:print0_s1_writedata -> print0:writedata
	wire         mm_interconnect_0_led_s1_chipselect;                       // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                         // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                          // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                            // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                        // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire         mm_interconnect_0_update_control_s1_chipselect;            // mm_interconnect_0:update_control_s1_chipselect -> update_control:chipselect
	wire  [31:0] mm_interconnect_0_update_control_s1_readdata;              // update_control:readdata -> mm_interconnect_0:update_control_s1_readdata
	wire   [1:0] mm_interconnect_0_update_control_s1_address;               // mm_interconnect_0:update_control_s1_address -> update_control:address
	wire         mm_interconnect_0_update_control_s1_write;                 // mm_interconnect_0:update_control_s1_write -> update_control:write_n
	wire  [31:0] mm_interconnect_0_update_control_s1_writedata;             // mm_interconnect_0:update_control_s1_writedata -> update_control:writedata
	wire         mm_interconnect_0_update_value_s1_chipselect;              // mm_interconnect_0:update_value_s1_chipselect -> update_value:chipselect
	wire  [31:0] mm_interconnect_0_update_value_s1_readdata;                // update_value:readdata -> mm_interconnect_0:update_value_s1_readdata
	wire   [1:0] mm_interconnect_0_update_value_s1_address;                 // mm_interconnect_0:update_value_s1_address -> update_value:address
	wire         mm_interconnect_0_update_value_s1_write;                   // mm_interconnect_0:update_value_s1_write -> update_value:write_n
	wire  [31:0] mm_interconnect_0_update_value_s1_writedata;               // mm_interconnect_0:update_value_s1_writedata -> update_value:writedata
	wire         mm_interconnect_0_x_coeff_bank_s1_chipselect;              // mm_interconnect_0:x_coeff_bank_s1_chipselect -> x_coeff_bank:chipselect
	wire  [31:0] mm_interconnect_0_x_coeff_bank_s1_readdata;                // x_coeff_bank:readdata -> mm_interconnect_0:x_coeff_bank_s1_readdata
	wire   [1:0] mm_interconnect_0_x_coeff_bank_s1_address;                 // mm_interconnect_0:x_coeff_bank_s1_address -> x_coeff_bank:address
	wire         mm_interconnect_0_x_coeff_bank_s1_write;                   // mm_interconnect_0:x_coeff_bank_s1_write -> x_coeff_bank:write_n
	wire  [31:0] mm_interconnect_0_x_coeff_bank_s1_writedata;               // mm_interconnect_0:x_coeff_bank_s1_writedata -> x_coeff_bank:writedata
	wire  [31:0] mm_interconnect_0_switch_s1_readdata;                      // switch:readdata -> mm_interconnect_0:switch_s1_readdata
	wire   [1:0] mm_interconnect_0_switch_s1_address;                       // mm_interconnect_0:switch_s1_address -> switch:address
	wire  [31:0] mm_interconnect_0_accel_yread_s1_readdata;                 // accel_yread:readdata -> mm_interconnect_0:accel_yread_s1_readdata
	wire   [1:0] mm_interconnect_0_accel_yread_s1_address;                  // mm_interconnect_0:accel_yread_s1_address -> accel_yread:address
	wire         mm_interconnect_0_y_coeff_bank_s1_chipselect;              // mm_interconnect_0:y_coeff_bank_s1_chipselect -> y_coeff_bank:chipselect
	wire  [31:0] mm_interconnect_0_y_coeff_bank_s1_readdata;                // y_coeff_bank:readdata -> mm_interconnect_0:y_coeff_bank_s1_readdata
	wire   [1:0] mm_interconnect_0_y_coeff_bank_s1_address;                 // mm_interconnect_0:y_coeff_bank_s1_address -> y_coeff_bank:address
	wire         mm_interconnect_0_y_coeff_bank_s1_write;                   // mm_interconnect_0:y_coeff_bank_s1_write -> y_coeff_bank:write_n
	wire  [31:0] mm_interconnect_0_y_coeff_bank_s1_writedata;               // mm_interconnect_0:y_coeff_bank_s1_writedata -> y_coeff_bank:writedata
	wire         mm_interconnect_0_print1_s1_chipselect;                    // mm_interconnect_0:print1_s1_chipselect -> print1:chipselect
	wire  [31:0] mm_interconnect_0_print1_s1_readdata;                      // print1:readdata -> mm_interconnect_0:print1_s1_readdata
	wire   [1:0] mm_interconnect_0_print1_s1_address;                       // mm_interconnect_0:print1_s1_address -> print1:address
	wire         mm_interconnect_0_print1_s1_write;                         // mm_interconnect_0:print1_s1_write -> print1:write_n
	wire  [31:0] mm_interconnect_0_print1_s1_writedata;                     // mm_interconnect_0:print1_s1_writedata -> print1:writedata
	wire  [31:0] mm_interconnect_0_accel_zread_s1_readdata;                 // accel_zread:readdata -> mm_interconnect_0:accel_zread_s1_readdata
	wire   [1:0] mm_interconnect_0_accel_zread_s1_address;                  // mm_interconnect_0:accel_zread_s1_address -> accel_zread:address
	wire         mm_interconnect_0_z_coeff_bank_s1_chipselect;              // mm_interconnect_0:z_coeff_bank_s1_chipselect -> z_coeff_bank:chipselect
	wire  [31:0] mm_interconnect_0_z_coeff_bank_s1_readdata;                // z_coeff_bank:readdata -> mm_interconnect_0:z_coeff_bank_s1_readdata
	wire   [1:0] mm_interconnect_0_z_coeff_bank_s1_address;                 // mm_interconnect_0:z_coeff_bank_s1_address -> z_coeff_bank:address
	wire         mm_interconnect_0_z_coeff_bank_s1_write;                   // mm_interconnect_0:z_coeff_bank_s1_write -> z_coeff_bank:write_n
	wire  [31:0] mm_interconnect_0_z_coeff_bank_s1_writedata;               // mm_interconnect_0:z_coeff_bank_s1_writedata -> z_coeff_bank:writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // accel_data_interrupt:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [accel_data_interrupt:reset_n, accel_xread:reset_n, accel_yread:reset_n, accel_zread:reset_n, cpu:reset_n, irq_mapper:reset, jtag_uart:rst_n, led:reset_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, print0:reset_n, print1:reset_n, rst_translator:in_reset, switch:reset_n, update_control:reset_n, update_value:reset_n, x_coeff_bank:reset_n, y_coeff_bank:reset_n, z_coeff_bank:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	nios2_cpu_accel_data_interrupt accel_data_interrupt (
		.clk        (clk_clk),                                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (mm_interconnect_0_accel_data_interrupt_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_accel_data_interrupt_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_accel_data_interrupt_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_accel_data_interrupt_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_accel_data_interrupt_s1_readdata),   //                    .readdata
		.in_port    (accel_interrupt_export),                               // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                              //                 irq.irq
	);

	nios2_cpu_accel_xread accel_xread (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_accel_xread_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_accel_xread_s1_readdata), //                    .readdata
		.in_port  (accel_xdata_export)                         // external_connection.export
	);

	nios2_cpu_accel_xread accel_yread (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_accel_yread_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_accel_yread_s1_readdata), //                    .readdata
		.in_port  (accel_ydata_export)                         // external_connection.export
	);

	nios2_cpu_accel_xread accel_zread (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_accel_zread_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_accel_zread_s1_readdata), //                    .readdata
		.in_port  (accel_zdata_export)                         // external_connection.export
	);

	nios2_cpu_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	nios2_cpu_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	nios2_cpu_led led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	nios2_cpu_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	nios2_cpu_print0 print0 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_print0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_print0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_print0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_print0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_print0_s1_readdata),   //                    .readdata
		.out_port   (disp0_export)                            // external_connection.export
	);

	nios2_cpu_print0 print1 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_print1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_print1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_print1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_print1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_print1_s1_readdata),   //                    .readdata
		.out_port   (disp1_export)                            // external_connection.export
	);

	nios2_cpu_switch switch (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_switch_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switch_s1_readdata), //                    .readdata
		.in_port  (switch_export)                         // external_connection.export
	);

	nios2_cpu_update_control update_control (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_update_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_update_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_update_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_update_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_update_control_s1_readdata),   //                    .readdata
		.out_port   (update_control_export)                           // external_connection.export
	);

	nios2_cpu_update_value update_value (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_update_value_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_update_value_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_update_value_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_update_value_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_update_value_s1_readdata),   //                    .readdata
		.out_port   (update_value_export)                           // external_connection.export
	);

	nios2_cpu_x_coeff_bank x_coeff_bank (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_x_coeff_bank_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_x_coeff_bank_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_x_coeff_bank_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_x_coeff_bank_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_x_coeff_bank_s1_readdata),   //                    .readdata
		.out_port   (x_coeff_bank_export)                           // external_connection.export
	);

	nios2_cpu_x_coeff_bank y_coeff_bank (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_y_coeff_bank_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_y_coeff_bank_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_y_coeff_bank_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_y_coeff_bank_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_y_coeff_bank_s1_readdata),   //                    .readdata
		.out_port   (y_coeff_bank_export)                           // external_connection.export
	);

	nios2_cpu_x_coeff_bank z_coeff_bank (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_z_coeff_bank_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_z_coeff_bank_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_z_coeff_bank_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_z_coeff_bank_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_z_coeff_bank_s1_readdata),   //                    .readdata
		.out_port   (z_coeff_bank_export)                           // external_connection.export
	);

	nios2_cpu_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                             (clk_clk),                                                   //                         clk_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                            // cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                 (cpu_data_master_address),                                   //                 cpu_data_master.address
		.cpu_data_master_waitrequest             (cpu_data_master_waitrequest),                               //                                .waitrequest
		.cpu_data_master_byteenable              (cpu_data_master_byteenable),                                //                                .byteenable
		.cpu_data_master_read                    (cpu_data_master_read),                                      //                                .read
		.cpu_data_master_readdata                (cpu_data_master_readdata),                                  //                                .readdata
		.cpu_data_master_write                   (cpu_data_master_write),                                     //                                .write
		.cpu_data_master_writedata               (cpu_data_master_writedata),                                 //                                .writedata
		.cpu_data_master_debugaccess             (cpu_data_master_debugaccess),                               //                                .debugaccess
		.cpu_instruction_master_address          (cpu_instruction_master_address),                            //          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest      (cpu_instruction_master_waitrequest),                        //                                .waitrequest
		.cpu_instruction_master_read             (cpu_instruction_master_read),                               //                                .read
		.cpu_instruction_master_readdata         (cpu_instruction_master_readdata),                           //                                .readdata
		.accel_data_interrupt_s1_address         (mm_interconnect_0_accel_data_interrupt_s1_address),         //         accel_data_interrupt_s1.address
		.accel_data_interrupt_s1_write           (mm_interconnect_0_accel_data_interrupt_s1_write),           //                                .write
		.accel_data_interrupt_s1_readdata        (mm_interconnect_0_accel_data_interrupt_s1_readdata),        //                                .readdata
		.accel_data_interrupt_s1_writedata       (mm_interconnect_0_accel_data_interrupt_s1_writedata),       //                                .writedata
		.accel_data_interrupt_s1_chipselect      (mm_interconnect_0_accel_data_interrupt_s1_chipselect),      //                                .chipselect
		.accel_xread_s1_address                  (mm_interconnect_0_accel_xread_s1_address),                  //                  accel_xread_s1.address
		.accel_xread_s1_readdata                 (mm_interconnect_0_accel_xread_s1_readdata),                 //                                .readdata
		.accel_yread_s1_address                  (mm_interconnect_0_accel_yread_s1_address),                  //                  accel_yread_s1.address
		.accel_yread_s1_readdata                 (mm_interconnect_0_accel_yread_s1_readdata),                 //                                .readdata
		.accel_zread_s1_address                  (mm_interconnect_0_accel_zread_s1_address),                  //                  accel_zread_s1.address
		.accel_zread_s1_readdata                 (mm_interconnect_0_accel_zread_s1_readdata),                 //                                .readdata
		.cpu_debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),             //             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                .write
		.cpu_debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                .read
		.cpu_debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                .readdata
		.cpu_debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                .writedata
		.cpu_debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                .byteenable
		.cpu_debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                .waitrequest
		.cpu_debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                .debugaccess
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                .chipselect
		.led_s1_address                          (mm_interconnect_0_led_s1_address),                          //                          led_s1.address
		.led_s1_write                            (mm_interconnect_0_led_s1_write),                            //                                .write
		.led_s1_readdata                         (mm_interconnect_0_led_s1_readdata),                         //                                .readdata
		.led_s1_writedata                        (mm_interconnect_0_led_s1_writedata),                        //                                .writedata
		.led_s1_chipselect                       (mm_interconnect_0_led_s1_chipselect),                       //                                .chipselect
		.onchip_memory2_0_s1_address             (mm_interconnect_0_onchip_memory2_0_s1_address),             //             onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write               (mm_interconnect_0_onchip_memory2_0_s1_write),               //                                .write
		.onchip_memory2_0_s1_readdata            (mm_interconnect_0_onchip_memory2_0_s1_readdata),            //                                .readdata
		.onchip_memory2_0_s1_writedata           (mm_interconnect_0_onchip_memory2_0_s1_writedata),           //                                .writedata
		.onchip_memory2_0_s1_byteenable          (mm_interconnect_0_onchip_memory2_0_s1_byteenable),          //                                .byteenable
		.onchip_memory2_0_s1_chipselect          (mm_interconnect_0_onchip_memory2_0_s1_chipselect),          //                                .chipselect
		.onchip_memory2_0_s1_clken               (mm_interconnect_0_onchip_memory2_0_s1_clken),               //                                .clken
		.print0_s1_address                       (mm_interconnect_0_print0_s1_address),                       //                       print0_s1.address
		.print0_s1_write                         (mm_interconnect_0_print0_s1_write),                         //                                .write
		.print0_s1_readdata                      (mm_interconnect_0_print0_s1_readdata),                      //                                .readdata
		.print0_s1_writedata                     (mm_interconnect_0_print0_s1_writedata),                     //                                .writedata
		.print0_s1_chipselect                    (mm_interconnect_0_print0_s1_chipselect),                    //                                .chipselect
		.print1_s1_address                       (mm_interconnect_0_print1_s1_address),                       //                       print1_s1.address
		.print1_s1_write                         (mm_interconnect_0_print1_s1_write),                         //                                .write
		.print1_s1_readdata                      (mm_interconnect_0_print1_s1_readdata),                      //                                .readdata
		.print1_s1_writedata                     (mm_interconnect_0_print1_s1_writedata),                     //                                .writedata
		.print1_s1_chipselect                    (mm_interconnect_0_print1_s1_chipselect),                    //                                .chipselect
		.switch_s1_address                       (mm_interconnect_0_switch_s1_address),                       //                       switch_s1.address
		.switch_s1_readdata                      (mm_interconnect_0_switch_s1_readdata),                      //                                .readdata
		.update_control_s1_address               (mm_interconnect_0_update_control_s1_address),               //               update_control_s1.address
		.update_control_s1_write                 (mm_interconnect_0_update_control_s1_write),                 //                                .write
		.update_control_s1_readdata              (mm_interconnect_0_update_control_s1_readdata),              //                                .readdata
		.update_control_s1_writedata             (mm_interconnect_0_update_control_s1_writedata),             //                                .writedata
		.update_control_s1_chipselect            (mm_interconnect_0_update_control_s1_chipselect),            //                                .chipselect
		.update_value_s1_address                 (mm_interconnect_0_update_value_s1_address),                 //                 update_value_s1.address
		.update_value_s1_write                   (mm_interconnect_0_update_value_s1_write),                   //                                .write
		.update_value_s1_readdata                (mm_interconnect_0_update_value_s1_readdata),                //                                .readdata
		.update_value_s1_writedata               (mm_interconnect_0_update_value_s1_writedata),               //                                .writedata
		.update_value_s1_chipselect              (mm_interconnect_0_update_value_s1_chipselect),              //                                .chipselect
		.x_coeff_bank_s1_address                 (mm_interconnect_0_x_coeff_bank_s1_address),                 //                 x_coeff_bank_s1.address
		.x_coeff_bank_s1_write                   (mm_interconnect_0_x_coeff_bank_s1_write),                   //                                .write
		.x_coeff_bank_s1_readdata                (mm_interconnect_0_x_coeff_bank_s1_readdata),                //                                .readdata
		.x_coeff_bank_s1_writedata               (mm_interconnect_0_x_coeff_bank_s1_writedata),               //                                .writedata
		.x_coeff_bank_s1_chipselect              (mm_interconnect_0_x_coeff_bank_s1_chipselect),              //                                .chipselect
		.y_coeff_bank_s1_address                 (mm_interconnect_0_y_coeff_bank_s1_address),                 //                 y_coeff_bank_s1.address
		.y_coeff_bank_s1_write                   (mm_interconnect_0_y_coeff_bank_s1_write),                   //                                .write
		.y_coeff_bank_s1_readdata                (mm_interconnect_0_y_coeff_bank_s1_readdata),                //                                .readdata
		.y_coeff_bank_s1_writedata               (mm_interconnect_0_y_coeff_bank_s1_writedata),               //                                .writedata
		.y_coeff_bank_s1_chipselect              (mm_interconnect_0_y_coeff_bank_s1_chipselect),              //                                .chipselect
		.z_coeff_bank_s1_address                 (mm_interconnect_0_z_coeff_bank_s1_address),                 //                 z_coeff_bank_s1.address
		.z_coeff_bank_s1_write                   (mm_interconnect_0_z_coeff_bank_s1_write),                   //                                .write
		.z_coeff_bank_s1_readdata                (mm_interconnect_0_z_coeff_bank_s1_readdata),                //                                .readdata
		.z_coeff_bank_s1_writedata               (mm_interconnect_0_z_coeff_bank_s1_writedata),               //                                .writedata
		.z_coeff_bank_s1_chipselect              (mm_interconnect_0_z_coeff_bank_s1_chipselect)               //                                .chipselect
	);

	nios2_cpu_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
